

 
 
 



 

window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /IF_Input_Table_tb/status
      waveform add -signals /IF_Input_Table_tb/IF_Input_Table_synth_inst/bmg_port/CLKA
      waveform add -signals /IF_Input_Table_tb/IF_Input_Table_synth_inst/bmg_port/ADDRA
      waveform add -signals /IF_Input_Table_tb/IF_Input_Table_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
